    Mac OS X            	   2  1     c                                      ATTR      c  �  �                 �     com.apple.lastuseddate#PS      �   *  $com.apple.metadata:_kMDItemUserTags       2  /com.apple.metadata:com_apple_mail_dateReceived     @   2  +com.apple.metadata:com_apple_mail_dateSent     r   *  5com.apple.metadata:com_apple_mail_isRemoteAttachment   �   �  %com.apple.metadata:kMDItemWhereFroms   M     com.apple.quarantine �]    ��3    bplist00�                            	bplist003A��ȸ                               bplist003A��ȱ                               bplist00                            	bplist00�_$Ilayda Yaman <ilaydayaman@gmail.com>VCNN tb_Pmessage:%3CCAHrs4Oy9i=5FH4_65QuF8AfoNNG5w4qg47e8DG26px1_BN24NQ@mail.gmail.com%3E3:                            �q/0082;5d975a16;Mail; 